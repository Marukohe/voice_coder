module fft_and_ifft();
    input clk;
    input [15:0] audio_in;

endmodule
