module mul_hanning();
endmodule;